bit strobe_tb;
mailbox#(int) mbx_tb = new();
event ev_tb;
